//
// Verilog Module CatRecognizer_lib.ControlUnit
//
// Created:
//          by - amitb.UNKNOWN (DESKTOP-GIFQ7HQ)
//          at - 16:06:27 17/11/2018
//
// using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
//

`resetall
`timescale 1ns/10ps
module ControlUnit ;


// ### Please start your Verilog code here ### 

endmodule
