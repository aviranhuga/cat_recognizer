library verilog;
use verilog.vl_types.all;
entity Neuron_tb is
end Neuron_tb;
